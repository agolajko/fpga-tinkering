/*
 * Copyright 2015 Forest Crossman
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *    http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 */

`include "cores/osdvu/uart.v"

module top(
	input iCE_CLK,
	input RS232_Rx_TTL,
	output RS232_Tx_TTL,
	output LED0,
	output LED1,
	output LED2,
	output LED3,
	output LED4,
    output PIO1_02,     // New output pin
    output PIO1_03,

	);

	wire reset = 0;
	reg transmit;
	reg [7:0] tx_byte;
	wire received;
	wire [7:0] rx_byte;
	wire is_receiving;
	wire is_transmitting;
	wire recv_error;

	assign LED4 = recv_error;

	uart #(
		.baud_rate(9600),                 // The baud rate in kilobits/s
		.sys_clk_freq(12000000)           // The master clock frequency
	)
	uart0(
		.clk(iCE_CLK),                    // The master clock for this module
		.rst(reset),                      // Synchronous reset
		.rx(RS232_Rx_TTL),                // Incoming serial line
		// .tx(RS232_Tx_TTL),                // Outgoing serial line
		.tx(PIO1_03),                // Outgoing serial line
		.transmit(transmit),              // Signal to transmit
		.tx_byte(tx_byte),                // Byte to transmit
		.received(received),              // Indicated that a byte has been received
		.rx_byte(rx_byte),                // Byte received
		.is_receiving(is_receiving),      // Low when receive line is idle
		.is_transmitting(is_transmitting),// Low when transmit line is idle
		.recv_error(recv_error)           // Indicates error in receiving packet.
	);


reg [24:0] counter = 0;  // Big enough counter to create visible delay


// assign LED0 = tx_byte; 
assign RS232_Tx_TTL = PIO1_03 ;  // Connect UART output to Pmod pin
assign LED0 = is_transmitting;
assign LED1 = is_transmitting;
assign LED2 = is_transmitting;
assign LED3 = is_transmitting;


always @(posedge iCE_CLK) begin
    counter <= counter + 1;
    
    if (counter == 0) begin  // Only transmit when counter rolls over
        tx_byte <= 8'b01010101;  // 0x55 = 'U'
        transmit <= 1;

	end


     else begin
        transmit <= 0;  // Need to drop transmit signal between sends

    end
end


endmodule
